
module struc_circuit_tb;

    reg a,b,c,d;
    wire y;


    struc_circuit(a,b,c,d,y);
    
    initial 
        begin
         
            a = 0;//1
            b = 0;
				c = 0;
				d = 0;
            #10; 
				
				a = 0;//2
            b = 0;
				c = 0;
				d = 1;
            #10; 
				
				a = 0;//3
            b = 0;
				c = 1;
				d = 0;
            #10; 
				
				a = 0;//4
            b = 0;
				c = 1;
				d = 1;
            #10;
				
				a = 0;//5
            b = 1;
				c = 0;
				d = 0;
            #10; 
				
				a = 0;//6
            b = 1;
				c = 0;
				d = 1;
            #10; 
				
				a = 0;//7
            b = 1;
				c = 1;
				d = 0;
            #10; 
				
				a = 0;//8
            b = 1;
				c = 1;
				d = 1;
            #10; 
				
				a = 1;//9
            b = 0;
				c = 0;
				d = 0;
            #10; 
				
				a = 1;//10
            b = 0;
				c = 0;
				d = 1;
            #10; 
				
				a = 1;//11
            b = 0;
				c = 1;
				d = 0;
            #10; 
				
				a = 1;//12
            b = 0;
				c = 1;
				d = 1;
            #10; 
				
				a = 1;//13
            b = 1;
				c = 0;
				d = 0;
            #10; 
				
				a = 1;//14
            b = 1;
				c = 0;
				d = 1;
            #10; 
				
				a = 1;//15
            b = 1;
				c = 1;
				d = 0;
            #10; 
				
				a = 1;//16
            b = 1;
				c = 1;
				d = 1;
            #10; 
						

           
endmodule