--test for VHDL code here
